library verilog;
use verilog.vl_types.all;
entity Mod_Teste_vlg_vec_tst is
end Mod_Teste_vlg_vec_tst;
